module show;
    initial begin
        $display("cc::::::::::::::::::;;:::;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;,,,,,,,,,,,,,,,,,,,,,,;;:oxkkOO00O0OOkOOo");
        $display("cc::::::::::::::::::::::;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;,,,,,,,,,,,,,,,,,,,,,,;;:lxkkOO00OOOOkO0o");
        $display("c:::::::::::::::::::::::::;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;,,,,,,,,,,,,,,,,,,,,,,;:lxkkkO00OOOOkO0d");
        $display("c::::::::::::::::::::::::;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;,,,,,,,,,,,,,,,,,,,,,,;:lxkkkO0OOOOOkO0d");
        $display("ccc::::::::::::::::::::;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;,,,,,,,,,,,,,,,,,,,,,,,;:lxkkkO00OOOOkO0x");
        $display("cc::::::::::::::::::::;;;;;;;;;;;;;;;;;;;:::ccccccccllllc:;;;;,,,,,,,,,,,,,,,,,,,,;:ldkkkO00OOOOkO0x");
        $display("c:::::::::::::::::::::::;;;;;;;;;;;;;:ldxOO0KXXXXXXNNNNXXKOxoc;,,,,,,,,,,,,,,,,,,,;;cdkkkO00OOOOkO0k");
        $display("::::::::::::::::::::::::;;;;;;;;;;;cdOKNNWWWWMMMMMMMMMMMMWWWNXOo:;;;,,,,,,,,,,,,,,;;cdkkkOOOOO0OO000");
        $display(":::::::::::::::::::::;;;;;;;;;;;;cokXWWWMMMMMMMMMMMMMMMMMMWWMWWXOo:;,;,,,,,,,,,,,,;;cdkkkOOOO0XXKKKK");  
        $display("c:::::::::::::::::::;;;;;;;;;:cldOXNWWMMMMMMMMMMMMMMMMMMMMMWWWWWWNOl;,,,,,,,,,,,,,;;cdkkkOO00XNNXXXX");
        $display("c:::::::::::::::::::;;;;;;:::ldkKWWWMMMMMMMMMMMMMMMMMMMMMMMMMWWWWWWXkc;,,,,,,,,,,,;;cdkkkOO0O0XXXXNX");
        $display("c::::::::::::::::::::;;;;;;::o0NWMMMMMMMMMMMMMMMMMMMMMMMMWWWMMMWWWWWN0l;,,,,,,,,,,,;:okkkkO0OkOO00XK");
        $display("cc:::::::::::::::::::;;;;;::lkNWWMMMMMMMMMMMMMMMMMMMMMMMMWWWWWWWWWWWWXx;,,,,,,,,,,,;:oxkkkO0OxkOkk00");
        $display(":c:::c::::::::::::::;;;;;::lkXWWWMMMMMMMMMMMMMMMMWWWWWWMMWWWNNNWNNWWNNOc;,,,,,,,,,,;:oxkkkO0OkkOOkO0");
        $display("cc::::::::::::::::::::::::cd0NWMMMMMMMMMMWWWMMMMWWWWNNNWWWWNNNNNNNNNNNKd;;,,,,,,,,,;:oxkkkO0OkOOOkk0");
        $display("ccc::c::::::::::::::::::::co0WWMMMMMMMMMMWWWWWNWWNNNNXXNNNNNXXXXNNNNNNNx:,,,,,,,,,,;:lxkkkOOOOOkkxk0");
        $display("cccccccc:::::::::::::::::::l0WMMMMMMMMWMMWWNXKKXXK000000000KXXXXXKXNNNNk:,,,,,,,,,,;:lxkkkOOOOOOkxk0");
        $display("ccccccccc::::::::::::::::::ckNMMMMWWWWWWWWNX0OkkOkxdllolldkOO0KNXkkKNWXx;,,,,,,,,,,;:lxkkkkO0OOOOkk0");
        $display("cccccccccc::::::::::::::::::oKWMWWWWWWNNNNNK00Okkkkkdolc::oxxxkXN0k0NWXo,,,,,,,,,,,;:lxkkkk00OOOOkk0");
        $display("ccccccccccccc:::::::::::::::ckNWWWWWWNXXXXK0Okxolclloolc:,,loox0XK00NW0c,,,,,,,,,,,;:lxkkkkO0OkOOkk0");
        $display("clccccccccccccc:::::::::::::cxKXWWWWNXK0Okxxkkkdoccc::;;,..;::cldxdkXNk:,,,,,,,,,,;;:lxkkkkO0OOOOkk0");
        $display("lllccccccccccccccc::::::::::lk0KXWWNXK0kdlccoxxddolcc:,,'..'';cddlldxkd;,,,,,,,,,,;;:ldkkkkO0OOOkkx0");
        $display("lllllllccccccccccccc::::::::cx00KNWNXK0koc;,,,;,,''''.'''.....',,',,,::,,,,,,,,,,,;;:ldkkkkO0OOOkkxO");
        $display("llllllllllcccccccccccccc:::::lO0KXNXXK0Odc;,''........',,'...........,,,,,,,,,,,,,;;:ldkkkkO00OOkkxk");
        $display("llllllllllllllllllcccccccccc:coOKKXKKK0Odl:,''.......';;;'...........',,,,,,,,,,,,;;:cdkkkkO00Okkkxk");
        $display("oooooloooooooooooooolllllllccccok00KKK0Oxl:;,'.......:ccl;..'.......'',,,,,,,,,,,,,;:cdkkkkO0Okkkkxk");
        $display("oooooooddddddddddddddooooooolllclkKXK00Oxoc;,'.......,;coc,,,.......',,,,,,,,,,,,,,;:cdkkkkO0Oxxkkxk");
        $display("dddxxxxxxxxxxxxddddddddddddooolllxXNXK0Oxoc:,''....................',,,,,,,,,,,,,,;;;cdxolokOOxxkkkk");
        $display("xxxxxxxxxxxxxxxxxxxxddddddddoooold0XKK0Oxoc:;,'.'''''',,,''''......',,,,,,,,,,,,,,,;;:oo,.'dOOkxkkkO");
        $display("kkkkkxxxxxxxxxxxxxxxxxxddddddooooodxOK0Okoc:;,,,,,,,:cllllcc:;,''.',,,,,,,,,,,,,,,;;;col,.,dOOkxkkxx");
        $display("kkkkkkkkkkkkkxxxxxxxxxxdddddddooooookKK0Oxl:;;,,,,,;:clc:;;;::,''',,,,,,,,,,,,,,,,,;;ldc,.,dOOO0K0Ok");
        $display("kkkkkkkkkkkkkkxxxxxxxxxxddddddooooookKK00kdl:;;;;;;;;;::::;;;,,,,,,,,,,,,,,,,,,,,,,;;lxl,.'lOOOKNXKK");
        $display("kkkkkkkkkkkkkkkxxxxxxxxxdddddddooood0K00OOkdoc:;;;;;;;,,,'''',,,,,,,,,,,,,,,,,,,,,,,;lxo;..:kOk0XNNN");
        $display("kkkkkkkkkkkkkkkkkxxxxxxxddddddddoooOKK0OOkkkxdlc:,,,,,,,,''''',,,,,,,,,,,,,,,,,,,,,,,cxo;..;dOkk0KXN");
        $display("OkkkOOOOkkkkkkkkkkxxxxxxxdddddddddkKK0Okkkkkxxddoc:;,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,;lxc'...ckkxkOKX");
        $display("OOOOOOOOOkkkkkkkkkxxxxxxxddddddodxO0Okddddxxxxxxxdoolcccccc;;,,,,,,,,,,,,,,,,,,,,,,,:dd,....,dkxkkO0");
        $display("OOOOOOOOkkkkkkkkkkkxxxxxdddddddddooxxdl:;:coddxxxxxddddool:;,,,,,,,,,,,,,,,,,,,,,,,,lxo,.....:oxkkkk");
        $display("OOOOOOOOkkkkkkkkkkkxxxxxxxxdoolc:;:cllc;'',;:cccllllllc:;;;;;;;;;;;;;;;;,,,,,,,,,,,;odc,'.....':dxxd");
        $display("OOOOOOkkkkkkkkkkkkkxxxxxddlc;,,''',;;:;'...'''''''''''''',;:;;;;;;;;;;;;,,,,,,,,,,,,,...........:odd");
        $display("OOOOOOOkkkkkkkkkkkkxxdolc;,'......'',''..................';:::;;,,''''''''',,,,,,;;..............:dd");
        $display("OkkOOOOOkkkkkkkkkxdolc;,,''..............................',;;:;;,''''''....'''''':c' ............,ld");
        $display("OOkOOOkkkkkkkkkkxoc::;,,''''.....''''''''''''''...........'';cc:,,''.............';;..............;l");
        $display("OOOOOOOkkkkkkkxdlc:;,''....................................',:llc;'''.......':c;..,;.  ...........',");
        $display("OOOOOOOOkkkxolc:,''...................    .................'',:lll:,'.......:O0Odcll'...''',,;,'...'");
        $display("OOOOOOOOkdl:;,''.....................        .................';cool:,......;k0000Oxlcclolc:;;'....'");
        $display("OOOOOOOxoc;,''.......    ......................................';coool:'.....:xO0Okxxddl:;'........,");
        $display("OOOOOOxoc;,'......         .....................................,codddoc;.....'oOOkxdol:;,,,,'''',,,");
        $display("OOOOOxo:;,'......            ...................................;ldddddol:'....,dOkxdlc::::::,,'',;,");
        $display("OO0Oxoc;,'......              ...............   ...............,codxdxdddol;'...,odol:,''',,;;,',;,'");
        $display("O00koc;,'.......            ..............       ............';codxxxxxxdddooc;,.':::::::clodooc:,'.");
        $display("O0Odl:;,'.........      ................             ......';codxxxxxxxxxxxxdddol:;;,''..';:lxxdl;..");
        $display("00koc;;,''..............................            .....,:lodxxxxxxxxxxxxxxxxxxddolc::;,,'.,oxdoc,.");
        $display("00xoc:;,,,'................'''..........          .....';coddxxxxxxxxxxxxxxxkkkkxxkkxxddoollldxddl:,");
        $display("\n\n\n");

            $display("                                               ..',,;:cccllc:;;,'..                                 ");
            $display("                                           ..,cokO00KKKKKKKK0000Okdoc;..                            ");
            $display("                                        .'cok0KKKKKKXKKKKXXXXKKKKKKKK0Od:..                         ");
            $display("                                      .cdOKKKKKKKKKKKKKKKXXXXXXXXXXXXK00Ox:.                        ");
            $display("                                    .ck0KKKKKKKKKKKKKKKKKKKKKKKKKXXXXXKKKK0x:..                     ");
            $display("                                  .;x0KKKKKKKKKKKKKKKKKK000OOO0000000KK00KXX0ko,.                   ");
            $display("                                 .cOKKKKKKKKKKKKKKKKKKK0kxoollllllllllllldx0XXK0o'                  ");
            $display("                                .cOKKKKKKKKKKKKKKKKKK0xl:,,'''',,,,'''',,;;ckXXXXk:.                ");
            $display("                               .;OKKKKKKKKKKKKKKKKKKko;'.................'',:dKXXXOc.               ");
            $display("                               'xKKKKKKKKKKKKKKKK0Oxc,'....................'':dKXXKO;               ");
            $display("                              .l000000KKKKKXKKK0koc:,''......................'ckKKK0o.              ");
            $display("                              ,x000000KKKKKK0kdl:,,,''........................;d0KKKx'              ");
            $display("                             .:O000000KKK0Oxlc:;,'''''...........  ...........,oO000d.              ");
            $display("                             .cO00000KKKOkdlc:;,,''''............   ..........'ck00Ol.              ");
            $display("                             .l000000K00kolc::::::;;,''......        .........'cO0Ox,               ");
            $display("                             .cO0O00K0K0kocc:cccc::;;,;;,'.....  .....'',,,,,''cOKOc.               ");
            $display("                              ,dkkkOKKK0kdollc:;'....'''''...........'......'''cOKd'                ");
            $display("                              .;llokKXKOdcccc:,'.',,:lc;,,',;;'..,,'';;;'',''',lkx;.                ");
            $display("                               ';:cdOK0koc:;,,'..''',;;'''':l:'.':;..,::'',,''':o;.                 ");
            $display("                               .;:coxOkdlc:;,''...........',;,...''...........':c.                  ");
            $display("                               .';::odoll:;,,'............''''.................''.                  ");
            $display("                                .',,:lllc:;,'.............','....................                   ");
            $display("                                 .',:llcc::;,...........,''''...................                    ");
            $display("                                  ,olccc::;;,'.........,;,'''..................                     ");
            $display("                                  ,Oklcc:;,,,'.........',,,,,,'................                     ");
            $display("                                  .:dl:::;,''.........''.......................                     ");
            $display("                                    .:c::;,'........,:;,,''''....'''''........                      ");
            $display("                                  ..cxocc:;,''......':c;,.........,c:'........                      ");
            $display("                                .'cdkkoclc:;,,'......';:;,'......','.........                       ");
            $display("                           ..',:lxkkOxc:lllc:;,''.....',;,''''..''.........                         ");
            $display("                      ...,:ldxxkkkkOko:,;cllcc:;,'..''...''''''...........                          ");
            $display("                  ..,;cldxxkkxxkkkkkko;,',;cccc::,,''................,;'...                         ");
            $display("             ..';:loddddxxxxxdxxkkkkxo;'.'',;:ccc:::;,'.............;cccc:;,'...                    ");
            $display("       ...';:cooddddddddddxxdddxxkxxdl;......',:::::::;;,'.........,clccccclllc:;,'...              ");
            $display("   ..';:lloooodooooooddddxxdddddxxxxdo:'........',;;;;;;;;;,''''...,llccccclllllcllcc:;'..          ");
            $display("  .coodddooddoddoooooddddxxdoodddxxxdo:'............',,,,''''...   .:lccclclllllllllllllc:,..       ");
            $display("  ,ddooddddoodoooooooooodxdooooddxxxdoc'........     ..',,'..      .,cccclllccllllllllllllll:,'..   ");
            $display("  ,odddoooooooooooooooooddoooooooddxdol,. .......      .''.         .:lclllclccllllllllllooolllc:.  ");
            $display("  ,oddddddddooooddooooodxdoooooolodxdooc.   .......   .';;,.        .:lcllllllllllllllllllloolooo,  ");
            $display("  ,oddddddoooooooooooooxxooooooooodddooo:.     .......::;:lc.       .;lcllllllllllllllllllloooooo,  ");
            $display("  ,odddddddooooooooooodxoloooooooooooooll,.     ....'okd:cdd;.      .;lllooollllllllllooooooooooo,  ");
            $display("  ,odoooooooooooooooodxdoooooooooooooooooc.     ....':xkoco:,'.     .;lllooollllllllloooooooooooo,  ");
            $display("  ,ddoodddoooodddooodxkxdoooollooooooodool;.   ......:xOdll,....    .,oollooolllooloooooooooddooo,  ");
            $display("  ,dddddddoodddddooooodxxxxoooooooooooooolc..   ....;x0kolc;. ...  ..,oooooooooooooodoooooddddddo,  ");
            $display("  ,odddddddoddododdddooodxkkdooooollooooool,..  ...;d00kolc:'. ......;ooooddooddodddddddddddddddo,  ");
            $display("  ,odddddddddddddddodddddxkxdoooolooooddooc;'.  .;ldO0Oxolcc:.   ....,ododddddddddddddddddddddxxd;  ");
            $display("  ;xddxddddddddddddddddxkxdoooodooooooddooo:,. .,dkkOOkolc:cl;.   ...;ddoddddddddddddxddddddddxxd;  ");
            $display("  ;xxdxxxddooddoddddddkkxdoooooddooooodddool:. .cxkOOOxoc::cll... ...,ddoddddddddddddxxdddxdxxxxd;  ");
            $display("  :kkxxkkxdooddddddddkOxddoodddoooooddddooooc'.,oxkOOkxoc::cll,. ....,ddddddxdddddddddxddxxxxxxxx;  ");
            $display("  :0K0OkkOxddddddddddk0Odoodddddddddddooooool'.:dxkOOkxolc:ccl;. ....;dxddddddddxxxxxxdxxxdxxxxxx;  ");
            $display("  ;k0KK0O00kxddddddddxOKkdoooodddddddddoddddl',ldxkkkkxdlccccl:. ....,dxddxxxddxxkkxxddxxxxkxxkkx:  ");
            $display("  ;kOO0KKKKKOxddddddxxk0Kkddddddddoooddoddddo;:oodxxxxxdlccc:c:......'oxdddxxxdxxxxkxxxxxxxxxxxkk:  ");
            $display("  ;xkkkOO0KXX0kxxddddxxkK0xdddddddddododddddoc:lodxxxxxolccc:c:'......lxddxxxxddxxxxxxxxxxxxkkxkk:  ");
            $display("  ;xkkkkkOOKNNKOkxddxxxxOKOxddddddddddddddddolllodddddddlccc:c:'......lxxdxxxxxdxxxxxxkxxxxxxxkOk:  ");
            $display("  :kkxxxxkkOKXNX0kxxddxxk0KOxdddddddddodddddddoloddddddolccccc:'......cxxxxxxxxxxxxxxxkxxxxxxkkOk:  ");
            $display("  cOOkxxxxxxkOKNX0kxxxxxxkKKkdddddddddooodddddoloooddddolllc::c,......ckkxxxxxxxxxxxxkkkxxxxxkkkx;  ");
            $display("  :0Okxxxxxddxxk0K0kdddxxxk0Oxdddoodddoooddddoollooooooolccc:::,.....'cxkddxxxxxxxxxxxxxxxxxxkkkx;  ");
            $display("\n\n\n");

            $display("kkkkxxkkxxkkkkkO000000KK0xddxxkO0Okkkkkkkkk0XXXXXXXXX0xddxxxxxxxoodoooooolooooooooolokOOOOOOOOOOOOOOOOOOO000OOOOOOOOOOOO");
            $display("xxxxdxxxxxxxxxk000000KXKxdxkOkxkxxxkkkxxxkk0KKKKXXXXKOxdxxxddddoloooooooolododddddoodkOkkOOOkOOOOOOOOOOOOOOOkkOOOOOOkkkk");
            $display("xdddddxxxxxxxxk0KK0KKKXOdoooolllcoxkkxxxxxk0KKKKKXXXKOxddxxddddoloddoooolllllllllllloxxxkkkkkkkkkkkkkkkkkkkkxxkkkkkkkkkk");
            $display("ddddddxxdddddxxk0KKKKKKkddxddxxdodxxxxxxxxk0KKKKXXXXX0OOO0Okkxdollllllllccllccccclccoxxxxxxxkkxxkkkxxxxxkkkxxxxxxxkkkkkx");
            $display("dxxxxddddddddddk0KKKKK0kdxkxddxdooxxxxddddk0KKXK00KKKXXXXXXXXXK0Oxolllcc:::;;:;;;::coxxxxxxxxxxxxxdddddxxxxxxxkkkkkkkkkk");
            $display("xkkOOxoodddddddk0KKKKK0kdxkxodxdlldddoooooxO0KOdoxkOOkOO00KKKKKXNXxcc::;,,'''',,,,,:odddddddddxddddddddxxxxxxkkkkkkkkkkk");
            $display("kkkOOoclddoodddk00KKKK0kodkxoodollooollllldOOxoclxOOxxk000000000K0xlc::;;;,,,,,,,,,:odddddddddddddooddddxxxdxxkkkkkkkkxx");
            $display("kkkOxc;collooooxO000000kodxdllooccccccccccdO0OkxooxxxkOO000O00Odcc:;,,,,'''''''''',cdddddooooddoooooddddxdddoddddxxxxxdd");
            $display("xxxxo,':ccllllldO000000xoodlcclc:;:::::::coOOOkxdooodxOO000000Odlcc:::;;;,,,,,,,,,;lodddolllllloooooooooddoooddddddddddd");
            $display("ddddl'.,:ccccllok000000xllclcc:::;;;:;;:::cllcccoxxxxkOkkOOOkkkkxxxddddoolcc:::;;,;loooolccccccllllllloooodooooooooooood");
            $display("olllc'.';:::ccclxOOOOOOxlccllc:,,;::;::c:::::;:clccloxxxdddddddddddoooodddddddddocclllollccclclllcclloooodddoooooooooooo");
            $display("llcc:...',;;;::cxOOOOOOdcc:cc:;'';lolc:,,,;;;:::ccllllcc:ccccclloooodoodxxddxxdddddoollccllllllllllloodddooooooodddddddd");
            $display("ccc::. .',,,;;;:dkkkkkkd:;,,::;,;:codo:,,;:cccccloolcc:;clcc::clloddddxkkxddoooooodolooooollcccllllooooooolllooooooddddd");
            $display("::::;. .''',,,,;okkkkkxl,,,:cc::loooxxoc::clllc:colc::;clllcccccldxdxxxO0kdoloooooollooddolccccccccccccllloooodooooooooo");
            $display(";:;;;. ...''',,;oxkkkkxo:,,,,;codxxkkxoc;:ccccccll:::::loollllcccloddxxkOOkdoooddxxdoollllccccccccccccccllloooooolllllll");
            $display(",;;;,.  ...'''',:ccccccc;,''',coxkO0kl;,;:ccccc::::;::clllllllllcclodxxkO00OxxxkO0Oo:ccccc::::::cccccccccllllllllllllooo");
            $display("'''''.........''...''''',,,,,;:ldxkOkc,,;:c:;;,,;:ccccclllllllllllllodxkO0kxxxkOOxocc:::c:::;;:ccllllllloooooooooooodddd");
            $display("...............'....''''''''',;:ldkOOd:::;;,,,,,;:cccllllllllllloolooddkOkddxkOxl:::::cccccc::cclllooooolloooooooooddddd");
            $display("........'''''''''....''''''',,,,;ldxOOxoc:;,,,,,,;:cclllllllllloooodddxxddxkkkdc;:cc::::::::ccllllclcccccllllllllllllooo");
            $display("'''''.....''',,,,,,,,,,,'''',,,,,;:ldxxkkxdolllclllllooodddddddddddddxxxxkkkdc:lxkkxl:::c::::ccccccc:::ccccccccclloooooo");
            $display("'''''''....''''''',,,,,;;,,,,,,,,'',:odxkO0KKXXKKKKKK0KKKKKKKK0OOOxdxxkOOO0kl;:d0KK0dccc:ccccccc:ccccccccccccccclloooddd");
            $display("........''''''''''''''''''''',,,,,,,,cdkO00KXXXXXXNNXKXXXNNNNNXK0kkkkO00KXX0o;:oxkkxl:cccc:::::::::cccclllcccccclllooddd");
            $display("...................................'',cx0KKKXKKXXNNNNXKKXXXNXNNXKKKXKXXNNNXOc,;;::::;;::::::::ccccccccccllllcccccclloool");
            $display(".......................................,lk0KKKXNNNNNNXKKKXXXNNXNNNNNNNNNNN0o;,;;::;;;;;:;;:::cccccccllllllccccccccccllll");
            $display("........................................,oOKKXXNNNNXXOk0KKXXXXXXNNNNNNNNNXx:,;;;;;;;,;;;;;::::::::ccccclllcccccccclloooo");
            $display("....................................''''';ldkO0000000dccdxkOOO0KXXXXXXXXKOo:;;;;;;;;;;;::::::::::::ccccccllllllllllooood");
            $display("...................'''''''''''''......'''',:oxkOOO00Oo,'',,;;;cdxkkOO0000kdlcccc::::;;;::::::::ccc::::cccllllccllllooooo");
            $display("''''''''''''''...'''''''''''''''''''''''''',cdkkOO0Ol,'''',,',;codddxkOO0Odcccloodddooolllcc:::::ccccccllllllllllllllllo");
            $display("'''''''''''''''''''''''''''''''''''',,,,,,,,;:clodxko;,,,,,,,,,;cooddkOO0xc;;;::ccllooddddddddoolllccccccllllllooooooooo");
            $display(",,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,;;:coxkO000000XKxlc::::::;::ccloxkOxl:::::c::::ccccloodddxxxxxxxxddddoooolllooooddd");
            $display(";;;;;;;;;;;;;;;;;,,;;;;;;;;;;;;;:coxkOO0KXNNNXXXKK00OOkxddoodooooc,,:oxkkdooooooooolooolloooooodddxxkkkOOOOOOkkkxxdddddd");
            $display(":::::;;;::::::::::::::::;;::::::cdkO00000OOkkxddooooooollllllllcok000KXNNK0OkxxxdddddddooooooooooooodddxxkkOOO0000000OOO");
            $display("llcccc::ccccc:ccccccc::c:::::::::::ccclcccccccc::ccccccccccccccccdOXXNNNNNNNXK0OkkxxxdddddddddddddddddoolooooddddxkkxkO0");
            $display("olllllllllclccccccclcccccccc:cccc:::::ccccccccccccccccclcclllllllld0XXXNNNNNNXK0Okxxdoooooooddooooooool:;:c:::c:;:c:;:dO");
            $display("\n\n\n");
    end

endmodule